LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE work.AluLib.all;

ENTITY Lab04 IS
END ENTITY;	

ARCHITECTURE q1 OF Lab04 IS
	SIGNAL a: INTEGER;
	SIGNAL b: INTEGER;
	SIGNAL op: BIT_VECTOR(1 DOWNTO 0);
	SIGNAL output: INTEGER;
BEGIN
	AluOutput: Alu PORT MAP(a,b,op,output);
END ARCHITECTURE;